module tlb();
  // TODO: associative memory

endmodule